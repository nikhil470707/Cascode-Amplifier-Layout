magic
tech scmos
timestamp 1731225671
<< nwell >>
rect 3 -3 42 37
rect 2 -61 41 -21
<< ntransistor >>
rect 12 -87 22 -85
rect 12 -120 22 -118
<< ptransistor >>
rect 10 17 34 19
rect 9 -41 33 -39
<< ndiffusion >>
rect 12 -77 22 -75
rect 12 -81 16 -77
rect 20 -81 22 -77
rect 12 -85 22 -81
rect 12 -91 22 -87
rect 12 -95 16 -91
rect 20 -95 22 -91
rect 12 -97 22 -95
rect 12 -110 22 -108
rect 12 -114 16 -110
rect 20 -114 22 -110
rect 12 -118 22 -114
rect 12 -124 22 -120
rect 12 -128 16 -124
rect 20 -128 22 -124
rect 12 -130 22 -128
<< pdiffusion >>
rect 10 28 34 31
rect 10 24 21 28
rect 25 24 34 28
rect 10 19 34 24
rect 10 12 34 17
rect 10 8 21 12
rect 25 8 34 12
rect 10 3 34 8
rect 9 -30 33 -27
rect 9 -34 20 -30
rect 24 -34 33 -30
rect 9 -39 33 -34
rect 9 -46 33 -41
rect 9 -50 20 -46
rect 24 -50 33 -46
rect 9 -55 33 -50
<< ndcontact >>
rect 16 -81 20 -77
rect 16 -95 20 -91
rect 16 -114 20 -110
rect 16 -128 20 -124
<< pdcontact >>
rect 21 24 25 28
rect 21 8 25 12
rect 20 -34 24 -30
rect 20 -50 24 -46
<< polysilicon >>
rect 1 17 10 19
rect 34 17 49 19
rect 0 -41 9 -39
rect 33 -41 48 -39
rect 10 -87 12 -85
rect 22 -87 25 -85
rect 10 -120 12 -118
rect 22 -120 25 -118
<< polycontact >>
rect -3 16 1 20
rect -4 -42 0 -38
rect 6 -88 10 -84
rect 6 -121 10 -117
<< metal1 >>
rect 25 24 46 28
rect -7 16 -3 20
rect 25 8 49 12
rect 46 -30 49 8
rect 24 -34 49 -30
rect -8 -42 -4 -38
rect 24 -50 48 -46
rect 45 -77 48 -50
rect 20 -81 48 -77
rect 2 -88 6 -84
rect 20 -95 48 -91
rect 44 -110 48 -95
rect 20 -114 48 -110
rect 2 -121 6 -117
rect 20 -128 26 -124
<< labels >>
rlabel metal1 45 25 45 25 7 vdd
rlabel metal1 -6 17 -6 17 3 vbias1
rlabel metal1 -6 -40 -6 -40 3 vbias2
rlabel metal1 3 -86 3 -86 1 vbias3
rlabel metal1 4 -119 4 -119 1 vin
rlabel metal1 24 -127 24 -127 1 gnd
rlabel metal1 47 -65 47 -65 7 vout
<< end >>
