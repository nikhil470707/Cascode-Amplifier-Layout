* Testbench for Cascode Amplifier
.INCLUDE "tsmc_spice_180nm.lib"
.INCLUDE "amp.spice"

* Voltage sources
VDD vdd 0 1.8
Vbias1 vbias1 0 1.12 ; 
Vbias2 vbias2 0 0.91
Vbias3 vbias3 0 0.87
Vin vin 0 SIN(0.6955 0.1 500k) ; 

* Simulation control
.TRAN 100p 10u ; 

.control
run
plot vin
plot vout
.endc

.end
