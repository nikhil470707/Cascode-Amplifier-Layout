magic
tech scmos
timestamp 1731222525
<< nwell >>
rect 531 145 570 187
rect 245 86 284 128
rect 324 86 363 128
rect 430 85 465 132
rect 528 87 567 129
<< ntransistor >>
rect 331 61 341 63
rect 432 63 442 65
rect 286 51 291 53
rect 485 63 495 65
rect 432 29 442 31
rect 485 29 495 31
rect 335 19 345 21
<< ptransistor >>
rect 539 165 563 167
rect 252 106 276 108
rect 332 106 356 108
rect 438 105 458 110
rect 536 107 560 109
<< ndiffusion >>
rect 331 72 341 75
rect 331 68 333 72
rect 337 68 341 72
rect 286 62 291 65
rect 290 58 291 62
rect 331 63 341 68
rect 432 73 442 77
rect 432 69 436 73
rect 440 69 442 73
rect 286 53 291 58
rect 331 57 341 61
rect 432 65 442 69
rect 485 73 495 77
rect 485 69 489 73
rect 493 69 495 73
rect 286 47 291 51
rect 331 53 333 57
rect 337 53 341 57
rect 331 49 341 53
rect 432 58 442 63
rect 485 65 495 69
rect 432 54 436 58
rect 440 54 442 58
rect 432 51 442 54
rect 485 58 495 63
rect 485 54 489 58
rect 493 54 495 58
rect 485 51 495 54
rect 290 43 291 47
rect 286 39 291 43
rect 432 39 442 43
rect 432 35 436 39
rect 440 35 442 39
rect 335 30 345 33
rect 335 26 337 30
rect 341 26 345 30
rect 432 31 442 35
rect 485 39 495 43
rect 485 35 489 39
rect 493 35 495 39
rect 335 21 345 26
rect 432 24 442 29
rect 485 31 495 35
rect 335 15 345 19
rect 432 20 436 24
rect 440 20 442 24
rect 432 17 442 20
rect 485 24 495 29
rect 485 20 489 24
rect 493 20 495 24
rect 485 17 495 20
rect 335 11 337 15
rect 341 11 345 15
rect 335 7 345 11
<< pdiffusion >>
rect 539 176 563 181
rect 539 172 548 176
rect 552 172 563 176
rect 539 167 563 172
rect 539 160 563 165
rect 539 156 548 160
rect 552 156 563 160
rect 539 151 563 156
rect 252 117 276 122
rect 252 113 263 117
rect 267 113 276 117
rect 252 108 276 113
rect 332 117 356 122
rect 332 113 341 117
rect 345 113 356 117
rect 252 101 276 106
rect 332 108 356 113
rect 438 121 458 126
rect 438 117 447 121
rect 451 117 458 121
rect 438 110 458 117
rect 536 118 560 123
rect 536 114 545 118
rect 549 114 560 118
rect 252 97 263 101
rect 267 97 276 101
rect 252 92 276 97
rect 332 101 356 106
rect 536 109 560 114
rect 332 97 341 101
rect 345 97 356 101
rect 332 92 356 97
rect 438 100 458 105
rect 438 96 447 100
rect 451 96 458 100
rect 438 91 458 96
rect 536 102 560 107
rect 536 98 545 102
rect 549 98 560 102
rect 536 93 560 98
<< ndcontact >>
rect 333 68 337 72
rect 286 58 290 62
rect 436 69 440 73
rect 489 69 493 73
rect 333 53 337 57
rect 436 54 440 58
rect 489 54 493 58
rect 286 43 290 47
rect 436 35 440 39
rect 337 26 341 30
rect 489 35 493 39
rect 436 20 440 24
rect 489 20 493 24
rect 337 11 341 15
<< pdcontact >>
rect 548 172 552 176
rect 548 156 552 160
rect 263 113 267 117
rect 341 113 345 117
rect 447 117 451 121
rect 545 114 549 118
rect 263 97 267 101
rect 341 97 345 101
rect 447 96 451 100
rect 545 98 549 102
<< polysilicon >>
rect 525 165 539 167
rect 563 165 573 167
rect 243 106 252 108
rect 276 106 290 108
rect 318 106 332 108
rect 356 106 366 108
rect 424 105 438 110
rect 458 105 467 110
rect 522 107 536 109
rect 560 107 570 109
rect 329 61 331 63
rect 341 61 343 63
rect 430 63 432 65
rect 442 63 444 65
rect 283 51 286 53
rect 291 51 293 53
rect 483 63 485 65
rect 495 63 498 65
rect 430 29 432 31
rect 442 29 444 31
rect 483 29 485 31
rect 495 29 498 31
rect 333 19 335 21
rect 345 19 347 21
<< polycontact >>
rect 521 164 525 168
rect 573 164 578 168
rect 239 105 243 109
rect 290 105 294 109
rect 314 105 318 109
rect 419 105 424 110
rect 467 105 472 110
rect 518 106 522 110
rect 325 60 329 64
rect 343 60 347 64
rect 426 62 430 66
rect 293 50 297 54
rect 444 62 448 66
rect 479 62 483 66
rect 426 28 430 32
rect 329 18 333 22
rect 444 28 448 32
rect 479 28 483 32
rect 347 18 351 22
<< metal1 >>
rect 482 176 527 177
rect 482 173 548 176
rect 482 147 489 173
rect 527 172 548 173
rect 520 164 521 168
rect 578 164 607 167
rect 573 163 607 164
rect 523 156 548 160
rect 523 148 528 156
rect 304 143 489 147
rect 520 143 528 148
rect 304 117 311 143
rect 421 121 427 143
rect 421 117 447 121
rect 520 118 525 143
rect 267 113 341 117
rect 520 114 545 118
rect 239 109 243 113
rect 294 105 314 109
rect 414 105 419 110
rect 472 106 518 110
rect 472 105 502 106
rect 267 97 293 101
rect 288 81 293 97
rect 316 97 341 101
rect 414 100 418 105
rect 316 83 321 97
rect 279 79 293 81
rect 318 82 321 83
rect 414 96 447 100
rect 520 98 545 102
rect 414 83 419 96
rect 520 90 525 98
rect 500 86 525 90
rect 500 83 508 86
rect 602 83 607 163
rect 318 79 363 82
rect 279 77 296 79
rect 279 76 297 77
rect 279 62 283 76
rect 293 64 297 76
rect 318 74 321 79
rect 414 79 449 83
rect 318 72 327 74
rect 444 73 449 79
rect 500 79 607 83
rect 500 74 505 79
rect 499 73 504 74
rect 318 70 333 72
rect 324 68 333 70
rect 440 69 449 73
rect 493 69 504 73
rect 420 64 426 66
rect 279 58 286 62
rect 293 60 325 64
rect 347 62 426 64
rect 448 62 479 66
rect 347 60 424 62
rect 293 54 297 60
rect 325 53 333 57
rect 440 54 451 58
rect 493 54 504 58
rect 280 43 286 47
rect 280 -15 284 43
rect 325 30 329 53
rect 446 39 451 54
rect 499 39 504 54
rect 440 35 451 39
rect 493 35 504 39
rect 325 26 337 30
rect 355 28 363 32
rect 373 28 426 32
rect 448 28 479 32
rect 355 22 359 28
rect 324 18 329 22
rect 351 18 359 22
rect 440 20 450 24
rect 493 20 504 24
rect 327 11 337 15
rect 327 -14 331 11
rect 446 -13 450 20
rect 500 -13 504 20
rect 446 -14 504 -13
rect 289 -15 504 -14
rect 280 -17 504 -15
rect 280 -18 450 -17
rect 280 -19 302 -18
rect 446 -20 450 -18
rect 500 -20 504 -17
<< m2contact >>
rect 363 77 373 82
rect 363 28 373 33
<< metal2 >>
rect 363 33 373 77
<< labels >>
rlabel metal1 444 22 444 22 1 gnd
rlabel metal1 428 119 428 119 1 Vdd
rlabel metal1 241 111 241 111 1 vbiasp
rlabel metal1 385 62 385 62 1 vbias3
rlabel metal1 387 29 387 29 1 vbias4
rlabel metal1 585 164 585 164 1 vbias1
rlabel metal1 512 108 512 108 1 vbias2
<< end >>
